module mul (
    input  [3:0] a,
    output reg [7:0] mul2,
    output reg [7:0] mul4,
    output reg [7:0] mul8,
    output reg       be4
);
    always @(*) begin
        /* */
    end
endmodule
