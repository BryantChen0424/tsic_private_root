module minmax (
    input  [7:0] a,
    input  [7:0] b,
    input        s,
    output reg [7:0] o
);
    always @(*) begin
        /* assignment */
    end
endmodule
