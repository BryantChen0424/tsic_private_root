module ops (
    input  [7:0] a,
    input  [7:0] b,
    input  [1:0] op,
    output reg [7:0] o,
    output reg overflow
);

    always @(*) begin

    end
endmodule
