module between (
    input  [7:0] a,
    output reg bt,
    output reg ubt
);
    always @(*) begin
        /* assignment */
    end
endmodule
